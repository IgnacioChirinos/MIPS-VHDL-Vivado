library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Instruction_Memory_IM is
	port (
		read_address: in STD_LOGIC_VECTOR (31 downto 0);
		instruction: out STD_LOGIC_VECTOR (31 downto 0)
	);
end Instruction_Memory_IM;

architecture Behavioral of Instruction_Memory_IM is

type memory is array (0 to 1023) of STD_LOGIC_VECTOR (7 downto 0);
signal Ins_Mem: memory := (


x"20",x"08",x"00",x"03",
x"20",x"09",x"00",x"03",
x"20",x"0A",x"00",x"03",
x"20",x"0B",x"00",x"03",
x"AC",x"08",x"00",x"24",
x"AC",x"09",x"00",x"28",
x"AC",x"0A",x"00",x"2C",
x"AC",x"0B",x"00",x"30",
x"20",x"19",x"00",x"02",
x"20",x"04",x"00",x"03",
x"20",x"05",x"00",x"02",
x"20",x"06",x"00",x"02",
x"20",x"07",x"00",x"03",
x"20",x"10",x"00",x"02",
x"20",x"11",x"00",x"02",
x"20",x"12",x"00",x"03",
x"20",x"13",x"00",x"02",
x"20",x"08",x"00",x"04",
x"20",x"09",x"00",x"01",
x"20",x"0A",x"00",x"03",
x"20",x"0B",x"00",x"02",
x"20",x"0C",x"00",x"02",
x"20",x"0D",x"00",x"02",
x"20",x"0E",x"00",x"03",
x"20",x"0F",x"00",x"03",
x"20",x"18",x"00",x"01",
x"8C",x"14",x"00",x"28",
x"8C",x"15",x"00",x"2C",
x"12",x"95",x"00",x"03",
x"20",x"10",x"00",x"01",
x"AC",x"10",x"00",x"34",
x"08",x"00",x"00",x"90",
x"03",x"28",x"A0",x"24",
x"00",x"C9",x"A8",x"24",
x"02",x"2A",x"B0",x"24",
x"02",x"95",x"A0",x"20",
x"02",x"96",x"A0",x"20",
x"AC",x"14",x"00",x"00",
x"00",x"88",x"A0",x"24",
x"00",x"E9",x"A8",x"24",
x"02",x"4A",x"B0",x"24",
x"02",x"95",x"A0",x"20",
x"02",x"96",x"A0",x"20",
x"AC",x"14",x"00",x"04",
x"00",x"A8",x"A0",x"24",
x"02",x"09",x"A8",x"24",
x"02",x"6A",x"B0",x"24",
x"02",x"95",x"A0",x"20",
x"02",x"96",x"A0",x"20",
x"AC",x"14",x"00",x"08",
x"03",x"2B",x"A0",x"24",
x"00",x"CC",x"A8",x"24",
x"02",x"2D",x"B0",x"24",
x"02",x"95",x"A0",x"20",
x"02",x"96",x"A0",x"20",
x"AC",x"14",x"00",x"0C",
x"00",x"8B",x"A0",x"24",
x"00",x"EC",x"A8",x"24",
x"02",x"4D",x"B0",x"24",
x"02",x"95",x"A0",x"20",
x"02",x"96",x"A0",x"20",
x"AC",x"14",x"00",x"10",
x"00",x"AB",x"A0",x"24",
x"02",x"0C",x"A8",x"24",
x"02",x"6D",x"B0",x"24",
x"02",x"95",x"A0",x"20",
x"02",x"96",x"A0",x"20",
x"AC",x"14",x"00",x"14",
x"03",x"2E",x"A0",x"24",
x"00",x"CF",x"A8",x"24",
x"02",x"38",x"B0",x"24",
x"02",x"95",x"A0",x"20",
x"02",x"96",x"A0",x"20",
x"AC",x"14",x"00",x"18",
x"00",x"8E",x"A0",x"24",
x"00",x"EF",x"A8",x"24",
x"02",x"58",x"B0",x"24",
x"02",x"95",x"A0",x"20",
x"02",x"96",x"A0",x"20",
x"AC",x"14",x"00",x"1C",
x"00",x"AE",x"A0",x"24",
x"02",x"0F",x"A8",x"24",
x"02",x"78",x"B0",x"24",
x"02",x"95",x"A0",x"20",
x"02",x"96",x"A0",x"20",
x"AC",x"14",x"00",x"20",
x"8C",x"08",x"00",x"00",
x"8C",x"09",x"00",x"04",
x"8C",x"0A",x"00",x"08",
x"8C",x"0B",x"00",x"0C",
x"8C",x"0C",x"00",x"10",
x"8C",x"0D",x"00",x"14",
x"8C",x"0E",x"00",x"18",
x"8C",x"0F",x"00",x"1C",
x"8C",x"18",x"00",x"20",
x"01",x"09",x"80",x"20",
x"02",x"0A",x"88",x"20",
x"02",x"2B",x"90",x"20",
x"02",x"4C",x"98",x"20",
x"02",x"6D",x"A0",x"20",
x"02",x"8E",x"A8",x"20",
x"02",x"AF",x"B0",x"20",
x"02",x"D8",x"B8",x"20",
x"12",x"E0",x"00",x"26",
x"8C",x"11",x"00",x"24",
x"8C",x"12",x"00",x"30",
x"12",x"32",x"00",x"01",
x"08",x"00",x"00",x"90",
x"20",x"10",x"00",x"02",
x"12",x"11",x"00",x"02",
x"20",x"10",x"00",x"03",
x"12",x"11",x"00",x"09",
x"20",x"10",x"00",x"01",
x"12",x"08",x"00",x"01",
x"08",x"00",x"00",x"90",
x"12",x"0C",x"00",x"01",
x"08",x"00",x"00",x"90",
x"10",x"09",x"00",x"01",
x"08",x"00",x"00",x"90",
x"10",x"0B",x"00",x"14",
x"08",x"00",x"00",x"90",
x"20",x"10",x"00",x"01",
x"12",x"08",x"00",x"01",
x"08",x"00",x"00",x"90",
x"12",x"0C",x"00",x"01",
x"08",x"00",x"00",x"90",
x"12",x"18",x"00",x"01",
x"08",x"00",x"00",x"90",
x"10",x"09",x"00",x"01",
x"08",x"00",x"00",x"90",
x"10",x"0A",x"00",x"01",
x"08",x"00",x"00",x"90",
x"10",x"0B",x"00",x"01",
x"08",x"00",x"00",x"90",
x"10",x"0D",x"00",x"01",
x"08",x"00",x"00",x"90",
x"10",x"0E",x"00",x"01",
x"08",x"00",x"00",x"90",
x"10",x"0F",x"00",x"01",
x"08",x"00",x"00",x"90",
x"AC",x"10",x"00",x"38",
x"08",x"00",x"00",x"90",
x"20",x"10",x"00",x"01",
x"AC",x"10",x"00",x"3C",
x"08",x"00",x"00",x"90",

--x"20",
--x"08",
--x"00",
--x"03",
--x"20",
--x"09",
--x"00",
--x"03",
--x"20",
--x"0A",
--x"00",
--x"03",
--x"20",
--x"0B",
--x"00",
--x"03",
--x"AC",
--x"08",
--x"00",
--x"24",
--x"AC",
--x"09",
--x"00",
--x"28",
--x"AC",
--x"0A",
--x"00",
--x"2c",
--x"AC",
--x"0B",
--x"00",
--x"30",
--x"20",
--x"08",
--x"00",
--x"02",
--x"20",
--x"09",
--x"00",
--x"03",
--x"20",
--x"0A",
--x"00",
--x"02",
--x"20",
--x"0B",
--x"00",
--x"02",
--x"20",
--x"0C",
--x"00",
--x"03",
--x"20",
--x"0D",
--x"00",
--x"02",
--x"20",
--x"0E",
--x"00",
--x"02",
--x"20",
--x"0F",
--x"00",
--x"03",
--x"20",
--x"18",
--x"00",
--x"02",
--x"AC",
--x"08",
--x"00",
--x"00",
--x"AC",
--x"09",
--x"00",
--x"04",
--x"AC",
--x"0A",
--x"00",
--x"08",
--x"AC",
--x"0B",
--x"00",
--x"0C",
--x"AC",
--x"0C",
--x"00",
--x"10",
--x"AC",
--x"0D",
--x"00",
--x"14",
--x"AC",
--x"0E",
--x"00",
--x"18",
--x"AC",
--x"0F",
--x"00",
--x"1C",
--x"AC",
--x"18",
--x"00",
--x"20",
--x"20",
--x"08",
--x"00",
--x"04",
--x"20",
--x"09",
--x"00",
--x"01",
--x"20",
--x"0A",
--x"00",
--x"03",
--x"20",
--x"0B",
--x"00",
--x"02",
--x"20",
--x"0C",
--x"00",
--x"02",
--x"20",
--x"0D",
--x"00",
--x"02",
--x"20",
--x"0E",
--x"00",
--x"03",
--x"20",
--x"0F",
--x"00",
--x"03",
--x"20",
--x"18",
--x"00",
--x"01",
--x"8C",
--x"10",
--x"00",
--x"28",
--x"8C",
--x"11",
--x"00",
--x"2c",
--x"12",
--x"11",
--x"00",
--x"03",
--x"20",
--x"12",
--x"00",
--x"01",
--x"AC",
--x"12",
--x"00",
--x"90",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"8C",
--x"10",
--x"00",
--x"00",
--x"8C",
--x"11",
--x"00",
--x"0C",
--x"8C",
--x"12",
--x"00",
--x"18",
--x"02",
--x"08",
--x"80",
--x"24",
--x"02",
--x"29",
--x"88",
--x"24",
--x"02",
--x"4A",
--x"90",
--x"24",
--x"02",
--x"11",
--x"98",
--x"20",
--x"02",
--x"72",
--x"A0",
--x"20",
--x"AC",
--x"14",
--x"00",
--x"34",
--x"8C",
--x"10",
--x"00",
--x"04",
--x"8C",
--x"11",
--x"00",
--x"10",
--x"8C",
--x"12",
--x"00",
--x"1C",
--x"02",
--x"08",
--x"80",
--x"24",
--x"02",
--x"29",
--x"88",
--x"24",
--x"02",
--x"4A",
--x"90",
--x"24",
--x"02",
--x"11",
--x"98",
--x"20",
--x"02",
--x"72",
--x"A0",
--x"20",
--x"AC",
--x"14",
--x"00",
--x"5C",
--x"38",
--x"10",
--x"00",
--x"08",
--x"8C",
--x"11",
--x"00",
--x"14",
--x"8C",
--x"12",
--x"00",
--x"20",
--x"02",
--x"08",
--x"80",
--x"24",
--x"02",
--x"29",
--x"88",
--x"24",
--x"02",
--x"4A",
--x"90",
--x"24",
--x"02",
--x"11",
--x"98",
--x"20",
--x"02",
--x"72",
--x"A0",
--x"20",
--x"AC",
--x"14",
--x"00",
--x"3c",
--x"8C",
--x"10",
--x"00",
--x"00",
--x"8C",
--x"11",
--x"00",
--x"0C",
--x"8C",
--x"12",
--x"00",
--x"18",
--x"02",
--x"0B",
--x"80",
--x"24",
--x"02",
--x"2C",
--x"88",
--x"24",
--x"02",
--x"4D",
--x"90",
--x"24",
--x"02",
--x"11",
--x"98",
--x"20",
--x"02",
--x"72",
--x"A0",
--x"20",
--x"AC",
--x"14",
--x"00",
--x"64",
--x"8C",
--x"10",
--x"00",
--x"04",
--x"8C",
--x"11",
--x"00",
--x"10",
--x"8C",
--x"12",
--x"00",
--x"1C",
--x"02",
--x"0B",
--x"80",
--x"24",
--x"02",
--x"2C",
--x"88",
--x"24",
--x"02",
--x"4D",
--x"90",
--x"24",
--x"02",
--x"11",
--x"98",
--x"20",
--x"02",
--x"72",
--x"A0",
--x"20",
--x"AC",
--x"14",
--x"00",
--x"68",
--x"8C",
--x"10",
--x"00",
--x"08",
--x"8C",
--x"11",
--x"00",
--x"14",
--x"8C",
--x"12",
--x"00",
--x"20",
--x"02",
--x"0B",
--x"80",
--x"24",
--x"02",
--x"2C",
--x"88",
--x"24",
--x"02",
--x"4D",
--x"90",
--x"24",
--x"02",
--x"11",
--x"98",
--x"20",
--x"02",
--x"72",
--x"A0",
--x"20",
--x"AC",
--x"14",
--x"00",
--x"6C",
--x"8C",
--x"10",
--x"00",
--x"00",
--x"8C",
--x"11",
--x"00",
--x"0C",
--x"8C",
--x"12",
--x"00",
--x"18",
--x"02",
--x"0E",
--x"80",
--x"24",
--x"02",
--x"2F",
--x"88",
--x"24",
--x"02",
--x"58",
--x"90",
--x"24",
--x"02",
--x"11",
--x"98",
--x"20",
--x"02",
--x"72",
--x"A0",
--x"20",
--x"AC",
--x"14",
--x"00",
--x"70",
--x"8C",
--x"10",
--x"00",
--x"04",
--x"8C",
--x"11",
--x"00",
--x"10",
--x"8C",
--x"12",
--x"00",
--x"1C",
--x"02",
--x"0E",
--x"80",
--x"24",
--x"02",
--x"2F",
--x"88",
--x"24",
--x"02",
--x"58",
--x"90",
--x"24",
--x"02",
--x"11",
--x"98",
--x"20",
--x"02",
--x"72",
--x"A0",
--x"20",
--x"AC",
--x"14",
--x"00",
--x"74",
--x"8C",
--x"10",
--x"00",
--x"08",
--x"8C",
--x"11",
--x"00",
--x"14",
--x"8C",
--x"12",
--x"00",
--x"20",
--x"02",
--x"0E",
--x"80",
--x"24",
--x"02",
--x"2F",
--x"88",
--x"24",
--x"02",
--x"58",
--x"90",
--x"24",
--x"02",
--x"11",
--x"98",
--x"20",
--x"02",
--x"72",
--x"A0",
--x"20",
--x"AC",
--x"14",
--x"00",
--x"78",
--x"8C",
--x"08",
--x"00",
--x"58",
--x"8C",
--x"09",
--x"00",
--x"5C",
--x"8C",
--x"0A",
--x"00",
--x"60",
--x"8C",
--x"0B",
--x"00",
--x"64",
--x"8C",
--x"0C",
--x"00",
--x"68",
--x"8C",
--x"0D",
--x"00",
--x"6C",
--x"8C",
--x"0E",
--x"00",
--x"70",
--x"8C",
--x"0F",
--x"00",
--x"74",
--x"8C",
--x"18",
--x"00",
--x"78",
--x"01",
--x"09",
--x"80",
--x"20",
--x"02",
--x"0A",
--x"88",
--x"20",
--x"02",
--x"2B",
--x"90",
--x"20",
--x"02",
--x"4C",
--x"98",
--x"20",
--x"02",
--x"6D",
--x"A0",
--x"20",
--x"02",
--x"8E",
--x"A8",
--x"20",
--x"02",
--x"AF",
--x"B0",
--x"20",
--x"02",
--x"D8",
--x"B8",
--x"20",
--x"12",
--x"C0",
--x"00",
--x"26",
--x"8C",
--x"11",
--x"00",
--x"48",
--x"8C",
--x"12",
--x"00",
--x"54",
--x"12",
--x"32",
--x"00",
--x"01",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"20",
--x"10",
--x"00",
--x"02",
--x"12",
--x"11",
--x"00",
--x"02",
--x"20",
--x"10",
--x"00",
--x"03",
--x"12",
--x"11",
--x"00",
--x"09",
--x"20",
--x"10",
--x"00",
--x"01",
--x"12",
--x"08",
--x"00",
--x"01",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"12",
--x"0C",
--x"00",
--x"01",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"10",
--x"09",
--x"00",
--x"01",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"10",
--x"0B",
--x"00",
--x"14",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"20",
--x"10",
--x"00",
--x"01",
--x"12",
--x"08",
--x"00",
--x"01",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"12",
--x"0C",
--x"00",
--x"01",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"12",
--x"18",
--x"00",
--x"01",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"10",
--x"09",
--x"00",
--x"01",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"10",
--x"0A",
--x"00",
--x"01",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"10",
--x"0B",
--x"00",
--x"01",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"10",
--x"0D",
--x"00",
--x"01",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"10",
--x"0E",
--x"00",
--x"01",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"10",
--x"0F",
--x"00",
--x"01",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"AC",
--x"10",
--x"00",
--x"7C",
--x"08",
--x"00",
--x"00",
--x"B4",
--x"20",
--x"10",
--x"00",
--x"01",
--x"AC",
--x"10",
--x"00",
--x"80",
--x"08",
--x"00",
--x"00",
--x"B4",
others => x"00"
);

begin	

--Instruction

instruction <= Ins_Mem(to_integer(unsigned(read_address)))&
               Ins_Mem(to_integer(unsigned(read_address))+1)&
               Ins_Mem(to_integer(unsigned(read_address))+2)&
               Ins_Mem(to_integer(unsigned(read_address))+3);
end Behavioral;